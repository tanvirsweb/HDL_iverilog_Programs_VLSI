module HalfAdder;
    initial begin
        $display("\nHello world,This is my 1st verilog program !!\n");
        $finish;
    end
endmodule

// D:\gitProjectsTanvirAnjomSiddique\000001HDL_Verilog\iverilog\bin\Verilog_Programs_HDL>iverilog -o 1 1.v       

// D:\gitProjectsTanvirAnjomSiddique\000001HDL_Verilog\iverilog\bin\Verilog_Programs_HDL>vvp 1   
// Hello world,This is my 1st verilog program !!
// 1.v:4: $finish called at 0 (1s)